`ifndef _FT_AsyncMode_vh_
`define _FT_AsyncMode_vh_
`include "../../hdl/FT_AsyncMode.v"
`endif //_FT_AsyncMode_vh_

`ifndef _FT_SyncMode_vh_
`define _FT_SyncMode_vh_
`include "../../hdl/FT_SyncMode.v"
`endif //_FT_SyncMode_vh_

`ifndef _dp_sync_fifo_vh_
`define _dp_sync_fifo_vh_
`include "../../hdl/dp_sync_fifo.v"
`endif //_dp_sync_fifo_vh_

`ifndef _FIFOlogicGated_vh_
`define _FIFOlogicGated_vh_
`include "../../hdl/FIFOlogicGated.v"
`endif //_FIFOlogicGated_vh_

`ifndef _dpram_vh_
`define _dpram_vh_
`include "../../hdl/dpram.v"
`endif //_dpram_vh_

`ifndef _FT2232_sim_vh_
`define _FT2232_sim_vh_
`include "../../hdl/FT2232_sim.v"
`endif //_FT2232_sim_vh_

`ifndef _spram_vh_
`define _spram_vh_
`include "../../hdl/spram.v"
`endif //_spram_vh_

`ifndef _FIFOlogicLUT_vh_
`define _FIFOlogicLUT_vh_
`include "../../hdl/FIFOlogicLUT.v"
`endif //_FIFOlogicLUT_vh_

`ifndef _sp_sync_fifo_vh_
`define _sp_sync_fifo_vh_
`include "../../hdl/sp_sync_fifo.v"
`endif //_sp_sync_fifo_vh_

`ifndef _dump_vh_
`define _dump_vh_
`include "../../include/dump.v"
`endif //_dump_vh_

